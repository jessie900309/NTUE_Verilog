module matrix8x8Rotate(clk,reset,segout,scanout);

input clk, reset;
output reg[7:0] segout;
output reg[2:0] scanout;
reg clk1;
reg [25:0] cnt_scan;
reg [25:0] clk_num = 12500000;
reg [7:0] q[0:7];

reg [2:0] Mode = 0; //000:start
reg [3:0] mode = 0;


//------------------ clock running -----------------------
	always@(posedge clk or negedge reset) begin
		if(!reset) begin
			cnt_scan<=0;
		end
		else begin
			cnt_scan<=cnt_scan+1;
			if(cnt_scan == clk_num) begin
				cnt_scan <=0;
				clk1 = ~clk1;
			end
		end
	end
//---------modify display digit ----------
	always @(posedge clk1, negedge reset) begin
		if (reset == 0) begin
			// reset matrix
			q[0] = 8'b11111111; q[1] = 8'b11111111; q[2] = 8'b11111111; q[3] = 8'b11111111;
			q[4] = 8'b11111111; q[5] = 8'b11111111; q[6] = 8'b11111111; q[7] = 8'b11111111;
			// reset mode&clock
			Mode <= 3'b000;
			mode <= 0;
			clk_num <= 12500000;
		end
		else begin
		
			case(Mode)
			
				3'b000://START
					if(mode==0)begin//S
						clk_num <= 12500000;
						q[0] = 8'b11100111;
						q[1] = 8'b11011011;
						q[2] = 8'b11011111;
						q[3] = 8'b11101111;
						q[4] = 8'b11110111;
						q[5] = 8'b11111011;
						q[6] = 8'b11011011;
						q[7] = 8'b11100111;
						mode <=1;
					end
					else if(mode==1)begin//T
						q[0] = 8'b11000001;
						q[1] = 8'b11110111;
						q[2] = 8'b11110111;
						q[3] = 8'b11110111;
						q[4] = 8'b11110111;
						q[5] = 8'b11110111;
						q[6] = 8'b11110111;
						q[7] = 8'b11110111;
						mode <=2;
					end
					else if(mode==2)begin//A
						q[0] = 8'b11100111;
						q[1] = 8'b11011011;
						q[2] = 8'b11011011;
						q[3] = 8'b11011011;
						q[4] = 8'b11000011;
						q[5] = 8'b11011011;
						q[6] = 8'b11011011;
						q[7] = 8'b11011011;
						mode <=3;
					end
					else if(mode==3)begin//R
						q[0] = 8'b10000111;
						q[1] = 8'b10111011;
						q[2] = 8'b10111011;
						q[3] = 8'b10000111;
						q[4] = 8'b10011111;
						q[5] = 8'b10101111;
						q[6] = 8'b10110111;
						q[7] = 8'b10111011;
						mode <=4;
					end
					else if(mode==4)begin//T
						q[0] = 8'b11000001;
						q[1] = 8'b11110111;
						q[2] = 8'b11110111;
						q[3] = 8'b11110111;
						q[4] = 8'b11110111;
						q[5] = 8'b11110111;
						q[6] = 8'b11110111;
						q[7] = 8'b11110111;
						Mode <= 3'b001;
						mode <=0;
					end
				
				3'b001: //fish slow
					if(mode==0)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=1;
					end
					else if(mode==1)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=2;
					end
					else if(mode==2)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=3;
					end
					else if(mode==3)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=4;
					end
					else if(mode==4)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						Mode <= 3'b010;
						mode <=0;
					end
				
				3'b010: //cat
					if(mode==0)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11101111;
						q[2] = 8'b11100111;
						q[3] = 8'b11000000;
						q[4] = 8'b10000000;
						q[5] = 8'b00000000;
						q[6] = 8'b00011000;
						q[7] = 8'b00011000;
						mode <=1;
					end
					else if(mode==1)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11110111;
						q[2] = 8'b11100111;
						q[3] = 8'b00000011;
						q[4] = 8'b00000001;
						q[5] = 8'b00000000;
						q[6] = 8'b00011000;
						q[7] = 8'b00011000;
						mode <=2;
					end
					else if(mode==2)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b01111110;
						q[2] = 8'b00111100;
						q[3] = 8'b00000000;
						q[4] = 8'b00000000;
						q[5] = 8'b00000000;
						q[6] = 8'b11000011;
						q[7] = 8'b11000011;
						Mode <= 3'b011;
						mode <=0;
					end
				
				3'b011: //fish fast
					if(mode==0)begin
						clk_num <= 1250000;
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=1;
					end
					else if(mode==1)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=2;
					end
					else if(mode==2)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=3;
					end
					else if(mode==3)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=4;
					end
					else if(mode==4)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=5;
					end
					else if(mode==5)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=6;
					end
					else if(mode==6)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=7;
					end
					else if(mode==7)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						mode <=8;
					end
					else if(mode==8)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b10001110;
						q[3] = 8'b01110100;
						q[4] = 8'b01111000;
						q[5] = 8'b10000100;
						q[6] = 8'b11111110;
						q[7] = 8'b11111111;
						mode <=9;
					end
					else if(mode==9)begin 
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111110;
						q[3] = 8'b10000100;
						q[4] = 8'b01111000;
						q[5] = 8'b01110100;
						q[6] = 8'b10001110;
						q[7] = 8'b11111111;
						Mode <= 3'b100;
						mode <=0;
					end
				
				3'b100: //fish dead
					if(mode==0)begin
						clk_num <= 50000000;
						q[0] = 8'b11100001;
						q[1] = 8'b11000011;
						q[2] = 8'b10000111;
						q[3] = 8'b10001111;
						q[4] = 8'b11011000;
						q[5] = 8'b01110100;
						q[6] = 8'b00001110;
						q[7] = 8'b10001111;
						Mode <=3'b111;
						mode <=0;
					end
				
				3'b111: //RIP
					if(mode==0) begin//R
						clk_num <= 25000000;
						q[0] = 8'b10000111;
						q[1] = 8'b10111011;
						q[2] = 8'b10111011;
						q[3] = 8'b10000111;
						q[4] = 8'b10011111;
						q[5] = 8'b10101111;
						q[6] = 8'b10110111;
						q[7] = 8'b10111011;
						mode <=1;
					end
					else if(mode==1) begin//I
						q[0] = 8'b11000001;
						q[1] = 8'b11110111;
						q[2] = 8'b11110111;
						q[3] = 8'b11110111;
						q[4] = 8'b11110111;
						q[5] = 8'b11110111;
						q[6] = 8'b11110111;
						q[7] = 8'b11000001;
						mode <=2;
					end
					else if(mode==2) begin//P
						q[0] = 8'b10000111;
						q[1] = 8'b10111011;
						q[2] = 8'b10111011;
						q[3] = 8'b10000111;
						q[4] = 8'b10111111;
						q[5] = 8'b10111111;
						q[6] = 8'b10111111;
						q[7] = 8'b10111111;
						mode <=3;
					end
					else if(mode==3) begin//end
						clk_num <= 75000000;
						q[0] = 8'b11111111;
						q[1] = 8'b01011010;
						q[2] = 8'b10111101;
						q[3] = 8'b01011010;
						q[4] = 8'b11111111;
						q[5] = 8'b11000011;
						q[6] = 8'b11000011;
						q[7] = 8'b11100111;
						mode <=4;
					end
					else if(mode==4) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b01011010;
						q[3] = 8'b10111101;
						q[4] = 8'b01011010;
						q[5] = 8'b11111111;
						q[6] = 8'b11000011;
						q[7] = 8'b11000011;
						mode <=5;
					end
					else if(mode==5) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b01011010;
						q[4] = 8'b10111101;
						q[5] = 8'b01011010;
						q[6] = 8'b11111111;
						q[7] = 8'b11000011;
						mode <=6;
					end
					else if(mode==6) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b11111111;
						q[4] = 8'b01011010;
						q[5] = 8'b10111101;
						q[6] = 8'b01011010;
						q[7] = 8'b11111111;
						mode <=7;
					end
					else if(mode==7) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b11111111;
						q[4] = 8'b11111111;
						q[5] = 8'b01011010;
						q[6] = 8'b10111101;
						q[7] = 8'b01011010;
						mode <=8;
					end
					else if(mode==8) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b11111111;
						q[4] = 8'b11111111;
						q[5] = 8'b11111111;
						q[6] = 8'b01011010;
						q[7] = 8'b10111101;
						mode <=9;
					end
					else if(mode==9) begin
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b11111111;
						q[4] = 8'b11111111;
						q[5] = 8'b11111111;
						q[6] = 8'b11111111;
						q[7] = 8'b01011010;
						mode <=10;
					end
					else if(mode==10) begin
						clk_num <= 125000000;
						q[0] = 8'b11111111;
						q[1] = 8'b11111111;
						q[2] = 8'b11111111;
						q[3] = 8'b11111111;
						q[4] = 8'b11111111;
						q[5] = 8'b11111111;
						q[6] = 8'b11111111;
						q[7] = 8'b11111111;
						Mode <=3'b000;
						mode <=0;
					end
			endcase
		end
	end
//-----------scan and display -------------
	always@(cnt_scan[15:13]) begin
		scanout <= cnt_scan[15:13];
	end
	
	always@(scanout) begin
		case(scanout)
			0: segout=q[0];
			1: segout=q[1];
			2: segout=q[2];
			3: segout=q[3];
			4: segout=q[4];
			5: segout=q[5];
			6: segout=q[6];
			7: segout=q[7];
			default: segout=8'b11111111;
		endcase 
	end
	
endmodule
